`include "uvm_macros.svh"
package fifo_pkg;
import uvm_pkg::*;
`include "transaction.sv"
`include "write_seq.sv"
`include "read_sequence.sv"
`include "write_sequencer.sv"
`include "read_sequencer.sv"
`include "virtual_sequencer.sv"
`include "virtual_sequence.sv"
`include "write_driver.sv"
`include "read_driver.sv"
`include "write_monitor.sv"
`include "read_monitor.sv"
`include "scoreboard.sv"
`include "subscriber.sv"
`include "write_agent.sv"
`include "read_agent.sv"
`include "environment.sv"
`include "test.sv"
endpackage
